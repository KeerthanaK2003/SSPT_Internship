module d_ff (
    input wire clk,
    input wire reset,
    input wire en,
    input wire d,
    output reg q
);

always @(posedge clk or posedge reset) begin
    if (reset)
        q <= 1'b0;
    else if (en)
        q <= d;
end

endmodule